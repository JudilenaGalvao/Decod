library verilog;
use verilog.vl_types.all;
entity Decod_vlg_vec_tst is
end Decod_vlg_vec_tst;
